module parser

import ast

fn (mut p Parser) top() {
}
