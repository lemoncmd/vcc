module parser

import (
  src2.ast
)

fn (p mut Parser) top() {
}
