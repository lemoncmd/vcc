module main

struct Type {
  kind []Typekind
}

enum Typekind {
  int
  pointer
}
