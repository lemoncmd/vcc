module parser

import ast

fn (p mut Parser) top() {
}
