module ast

struct ScopeTable {}

